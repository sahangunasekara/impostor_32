`timescale 1ns/100ps

module load(input clk, input [31:0] pc_out, input reset, output [31:0] ALU_result);

	//PC pc (.clk(clk), .reset(rst))
	
  wire [31:0] instruction,ScrB;
	wire [1:0] Alu_op;
	wire [3:0] out_to_alu;
   wire [1:0] equal_comp;
	wire [2:0] mem;
	wire RegWrite, MemWrite, MemRead, Branch, ALUSrc,jump, ALU_En, mem_reg,zero;
	
	wire [4:0] read_addr_1; 
	wire [4:0] read_addr_2; 
	wire [4:0] write_addr;
	wire [31:0] write_data;
	wire [31:0] read_data_1;
	wire [31:0] read_data_2;
	wire [6:0] Opcode;
	wire [31:0] immidiate;
	wire [3:0] funct;
	wire [31:0] read_data;

	
	
	//wire reg_w;
instruction_memory Instruction_memory (
	.read_addr(pc_out), 
	.clk(clk), 
	.instruction(instruction)
	);
	
mux_N_bit #(32) data_memory_mux (
		.in0(ALU_result), 
		.in1(read_data), 
		.mux_out(write_data), 
		.control(mem_reg)
		);

instruction_parser instruction_parser(
		.instruction(instruction),
		.rs1(read_addr_1),
		.rs2(read_addr_2),
		.rd(write_addr),
		.opcode(Opcode),
		.imm(immidiate),
		.func(funct)
		);
	
	// for R type instruction
register_file register_file(
    .clk(clk),
    .read_addr_1(read_addr_1),
    .read_addr_2(read_addr_2),
    .write_addr(write_addr),
    .write_data(write_data),//..........
    .reg_write(RegW),
  	 .read_data_1(read_data_1),
    .read_data_2(read_data_2)
	 );
	
alu_control ALU_control (
	.funct(funct),
	.alu_op(Alu_op),
	.out_to_alu(out_to_alu),
	.ALU_En(ALU_En),
	.equal_comp(equal_comp),
	.mem(mem)
 
	);
maincontroller contr(
	.Opcode(Opcode),
	.RegWrite(RegW), 
	.MemWrite(MemW), 
	.MemRead(MemR), 
	.Branch(Branch), 
	.ALUSrc( ALUSrc), 
	.Aluop(Alu_op),
	.jump(jump), 
	.ALU_En(ALU_En), 
	.mem_reg(mem_reg)
	);
	
data_memory data_memory_module(
    .clk(clk),
    .mem_read(MemR),
    .mem_write(MemW),
    .DATA_MEM_In(mem),
    .read_data(read_data),
    .write_data(read_data_2),
    .addr(ALU_result)
    // Add other inputs and outputs here
  );
  
mux_N_bit #(32) ALU_mux (
		.in0(read_data_2), 
		.in1(immidiate), 
		.mux_out(ScrB), 
		.control(  ALUSrc)
		);	
alu sahan(
  	.ScrA(read_data_1),
  	.ScrB(ScrB),
	.alu_control(out_to_alu),
	.ALUResult(ALU_result),
	.zero(zero),
	.equalComp(equal_comp)
	);
endmodule